netcdf soildata {
dimensions:
  lon = xlen ;
  lat = ylen ;
  depth = 6 ;
  nb = 2 ;

variables:

  double lon(lon) ;
    lon:long_name = "longitude" ;
    lon:units = "degrees_east" ;
    lon:actual_range = 0., 0. ;
    lon:axis = "X" ;

  double lat(lat) ;
    lat:long_name = "latitude" ;
    lat:units = "degrees_north" ;
    lat:actual_range = 0., 0. ;
    lat:axis = "Y" ;

  float depth(depth) ;
    depth:long_name = "vertical position of layer midpoint (below soil surface)" ;
    depth:units = "cm" ;
    depth:positive = "down" ;
    depth:bounds = "layer_bnds" ;
    depth:axis = "Z" ;
    
  float layer_bnds(depth,nb) ;
    layer_bnds:units = "cm" ;
    layer_bnds:positive = "down" ;

  float dz(depth) ;
    dz:long_name = "soil layer thickness" ;
    dz:units = "cm" ;

  byte WRB(lat, lon) ;
    WRB:long_name = "Predicted WRB 2006 subgroup classes" ;
    WRB:units = "class" ;
    WRB:_FillValue = -1b ;
    WRB:missing_value = -1b ;
    WRB:actual_range = 0b, -1b ;
    WRB:valid_range = 1b, 118b ;
    WRB:source = "SoilGrids 2017" ;
    WRB:_Storage = "chunked" ;
    WRB:_ChunkSizes = ylen, xlen ;
    WRB:_DeflateLevel = 1 ;

  byte USDA(lat, lon) ;
    USDA:long_name = "Predicted USDA 2014 suborder classes" ;
    USDA:units = "class" ;
    USDA:_FillValue = -1b ;
    USDA:missing_value = -1b ;
    USDA:actual_range = 0b, -1b ;
    USDA:valid_range = 1b, 99b ;
    USDA:source = "SoilGrids 2017" ;
    USDA:_Storage = "chunked" ;
    USDA:_ChunkSizes = ylen, xlen ;
    USDA:_DeflateLevel = 1 ;

  float thickness(lat, lon) ;
    thickness:long_name = "average soil and sedimentary deposit thickness" ;
    thickness:units = "m" ;
    thickness:_FillValue = -9999.f ;
    thickness:missing_value = -9999.f ;
    thickness:actual_range = 100.f, -100.f ;
    thickness:source = "Pelletier et al., 2016" ;
    thickness:_Storage = "chunked" ;
    thickness:_ChunkSizes = ylen, xlen ;
    thickness:_DeflateLevel = 1 ;
    
  short sand(depth, lat, lon) ;
    sand:long_name = "sand content by mass" ;
    sand:units = "fraction" ;
    sand:_FillValue = -32768s ;
    sand:missing_value = -32768s ;
    sand:actual_range = 100.f, -100.f ;
    sand:valid_range = 0s, 1000s ;
    sand:scale_factor = 0.001f ;
    sand:source = "SoilGrids 2020" ;
    sand:_Storage = "chunked" ;
    sand:_Shuffle = "true" ;
    sand:_ChunkSizes = 1, ylen, xlen ;
    sand:_DeflateLevel = 1 ;

  short silt(depth, lat, lon) ;
    silt:long_name = "silt content by mass" ;
    silt:units = "fraction" ;
    silt:_FillValue = -32768s ;
    silt:missing_value = -32768s ;
    silt:actual_range = 100.f, -100.f ;
    silt:valid_range = 0s, 1000s ;
    silt:scale_factor = 0.001f ;
    silt:source = "SoilGrids 2020" ;
    silt:_Storage = "chunked" ;
    silt:_Shuffle = "true" ;
    silt:_ChunkSizes = 1, ylen, xlen ;
    silt:_DeflateLevel = 1 ;

  short clay(depth, lat, lon) ;
    clay:long_name = "clay content by mass" ;
    clay:units = "fraction" ;
    clay:_FillValue = -32768s ;
    clay:missing_value = -32768s ;
    clay:actual_range = 100.f, -100.f ;
    clay:valid_range = 0s, 1000s ;
    clay:scale_factor = 0.001f ;
    clay:source = "SoilGrids 2020" ;
    clay:_Storage = "chunked" ;
    clay:_Shuffle = "true" ;
    clay:_ChunkSizes = 1, ylen, xlen ;
    clay:_DeflateLevel = 1 ;

  short cfvo(depth, lat, lon) ;
    cfvo:long_name = "coarse fragments by volume" ;
    cfvo:units = "fraction" ;
    cfvo:_FillValue = -32768s ;
    cfvo:missing_value = -32768s ;
    cfvo:actual_range = 100.f, -100.f ;
    cfvo:valid_range = 0s, 1000s ;
    cfvo:scale_factor = 0.001f ;
    cfvo:source = "SoilGrids 2020" ;
    cfvo:_Storage = "chunked" ;
    cfvo:_Shuffle = "true" ;
    cfvo:_ChunkSizes = 1, ylen, xlen ;
    cfvo:_DeflateLevel = 1 ;

  short soc(depth, lat, lon) ;
    soc:long_name = "Soil organic carbon content by mass" ;
    soc:units = "fraction" ;
    soc:_FillValue = -32768s ;
    soc:missing_value = -32768s ;
    soc:actual_range = 100.f, -100.f ;
    soc:valid_range = 0s, 10000s ;
    soc:scale_factor = 0.0001f ;
    soc:source = "SoilGrids 2020" ;
    soc:_Storage = "chunked" ;
    soc:_Shuffle = "true" ;
    soc:_ChunkSizes = 1, ylen, xlen ;
    soc:_DeflateLevel = 1 ;

  short bdod(depth, lat, lon) ;
    bdod:long_name = "SoilGrids bulk density" ;
    bdod:units = "g cm-3" ;
    bdod:_FillValue = -32768s ;
    bdod:missing_value = -32768s ;
    bdod:actual_range = 0.f, 0.f ;
    bdod:scale_factor = 0.01f ;
    bdod:source = "SoilGrids 2020" ;
    bdod:_Storage = "chunked" ;
    bdod:_ChunkSizes = 1, ylen, xlen ;
    bdod:_DeflateLevel = 1 ;

  float bulk(depth, lat, lon) ;
    bulk:long_name = "calculated bulk density" ;
    bulk:units = "g cm-3" ;
    bulk:_FillValue = -9999.f ;
    bulk:missing_value = -9999.f ;
    bulk:actual_range = 100.f, -100.f ;
    bulk:source = "Balland et al., 2008" ;
    bulk:_Storage = "chunked" ;
    bulk:_ChunkSizes = 1, ylen, xlen ;
    bulk:_DeflateLevel = 1 ;

  float Tsat(depth, lat, lon) ;
    Tsat:long_name = "soil porosity (Theta-sat)" ;
    Tsat:units = "fraction" ;
    Tsat:_FillValue = -9999.f ;
    Tsat:missing_value = -9999.f ;
    Tsat:actual_range = 100.f, -100.f ;
    Tsat:source = "Sandoval et al., 2024" ;
    Tsat:_Storage = "chunked" ;
    Tsat:_ChunkSizes = 1, ylen, xlen ;
    Tsat:_DeflateLevel = 1 ;

  float T33(depth, lat, lon) ;
    T33:long_name = "soil water content at field capacity (-33 kPa)" ;
    T33:units = "mm cm-1" ;
    T33:_FillValue = -9999.f ;
    T33:missing_value = -9999.f ;
    T33:actual_range = 100.f, -100.f ;
    T33:source = "Sandoval et al., 2024" ;
    T33:_Storage = "chunked" ;
    T33:_ChunkSizes = 1, ylen, xlen ;
    T33:_DeflateLevel = 1 ;

  float T1500(depth, lat, lon) ;
    T1500:long_name = "soil water content at permanent wilting point (-1500 kPa)" ;
    T1500:units = "mm cm-1" ;
    T1500:_FillValue = -9999.f ;
    T1500:missing_value = -9999.f ;
    T1500:actual_range = 100.f, -100.f ;
    T1500:source = "Sandoval et al., 2024" ;
    T1500:_Storage = "chunked" ;
    T1500:_ChunkSizes = 1, ylen, xlen ;
    T1500:_DeflateLevel = 1 ;

  float whc(depth, lat, lon) ;
    whc:long_name = "water holding capacity defined as T33-T1500, reduced for coarse fragment volume" ;
    whc:units = "mm cm-1" ;
    whc:_FillValue = -9999.f ;
    whc:missing_value = -9999.f ;
    whc:actual_range = 100.f, -100.f ;
    whc:_Storage = "chunked" ;
    whc:_ChunkSizes = 1, ylen, xlen ;
    whc:_DeflateLevel = 1 ;

  float Ksat(depth, lat, lon) ;
    Ksat:long_name = "saturated hydraulic conductivity" ;
    Ksat:units = "mm h-1" ;
    Ksat:_FillValue = -9999.f ;
    Ksat:missing_value = -9999.f ;
    Ksat:actual_range = 100.f, -100.f ;
    Ksat:source = "Sandoval et al., 2024 (code only)" ;
    Ksat:_Storage = "chunked" ;
    Ksat:_ChunkSizes = 1, ylen, xlen ;

// global attributes:
    :Conventions = "CF-1.11" ;
    :title = "Primary and derived soil properties" ;
    :citation1 = "Hengl, T., Mendes de Jesus, J., Heuvelink, G. B., Ruiperez Gonzalez, M., Kilibarda, M., Blagotic, A., Shangguan, W., Wright, M. N., Geng, X., Bauer-Marschallinger, B., Guevara, M. A., Vargas, R., MacMillan, R. A., Batjes, N. H., Leenaars, J. G., Ribeiro, E., Wheeler, I., Mantel, S., & Kempen, B. (2017). SoilGrids250m: Global gridded soil information based on machine learning. PLoS One, 12(2), e0169748. doi:10.1371/journal.pone.0169748" ;
    :citation2 = "Pelletier, J. D., Broxton, P. D., Hazenberg, P., Zeng, X., Troch, P. A., Niu, G. Y., Williams, Z., Brunke, M. A., & Gochis, D. (2016). A gridded global data set of soil, intact regolith, and sedimentary deposit thicknesses for regional and global land surface modeling. Journal of Advances in Modeling Earth Systems, 8(1), 41-65. doi:10.1002/2015ms000526" ;
    :citation4 = "Balland, V., Pollacco, J. A. P., & Arp, P. A. (2008). Modeling soil hydraulic properties for a wide range of soil conditions. Ecological Modelling, 219(3-4), 300-316. doi:10.1016/j.ecolmodel.2008.07.009" ;
    :citation3 = "Sandoval, D., Prentice, I. C., & Nóbrega, R. L. B. (2024). Simple process-led algorithms for simulating habitats (SPLASH v.2.0): robust calculations of water and energy fluxes. Geoscientific Model Development, 17(10), 4229-4309. doi:10.5194/gmd-17-4229-2024" ;
    :node_offset = 1 ;

}
