netcdf soildata {
dimensions:
	lon = xlen ;
	lat = ylen ;
	depth = 6 ;
	nb = 2 ;

variables:

	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:actual_range = 0., 0. ;
		lon:axis = "X" ;

	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:actual_range = 0., 0. ;
		lat:axis = "Y" ;

	float depth(depth) ;
		depth:long_name = "depth_below_land" ;
		depth:units = "cm" ;
		depth:positive = "down" ;
		depth:bounds = "layer_bnds" ;
		depth:axis = "Z" ;
		
	float layer_bnds(depth,nb) ;
		layer_bnds:units = "cm" ;
		layer_bnds:positive = "down" ;

	float dz(depth) ;
		dz:long_name = "soil layer thickness" ;
		dz:units = "cm" ;

	byte soiltype(lat, lon) ;
		soiltype:long_name = "Predicted WRB 2006 subgroup" ;
		soiltype:units = "class" ;
		soiltype:_FillValue = -1b ;
		soiltype:missing_value = -1b ;
		soiltype:actual_range = 0b, -1b ;
		soiltype:valid_range = 1b, 118b ;
		soiltype:_Storage = "chunked" ;
		soiltype:_ChunkSizes = ylen, xlen ;
		soiltype:_DeflateLevel = 1 ;

	short sand(depth, lat, lon) ;
		sand:long_name = "sand content by mass" ;
		sand:units = "fraction" ;
		sand:_FillValue = -32768s ;
		sand:missing_value = -32768s ;
		sand:actual_range = 100.f, -100.f ;
		sand:valid_range = 0s, 1000s ;
		sand:scale_factor = 0.001f ;
		sand:_Storage = "chunked" ;
		sand:_Shuffle = "true" ;
		sand:_ChunkSizes = 1, ylen, xlen ;
		sand:_DeflateLevel = 1 ;

	short silt(depth, lat, lon) ;
		silt:long_name = "silt content by mass" ;
		silt:units = "fraction" ;
		silt:_FillValue = -32768s ;
		silt:missing_value = -32768s ;
		silt:actual_range = 100.f, -100.f ;
		silt:valid_range = 0s, 1000s ;
		silt:scale_factor = 0.001f ;
		silt:_Storage = "chunked" ;
		silt:_Shuffle = "true" ;
		silt:_ChunkSizes = 1, ylen, xlen ;
		silt:_DeflateLevel = 1 ;

	short clay(depth, lat, lon) ;
		clay:long_name = "clay content by mass" ;
		clay:units = "fraction" ;
		clay:_FillValue = -32768s ;
		clay:missing_value = -32768s ;
		clay:actual_range = 100.f, -100.f ;
		clay:valid_range = 0s, 1000s ;
		clay:scale_factor = 0.001f ;
		clay:_Storage = "chunked" ;
		clay:_Shuffle = "true" ;
		clay:_ChunkSizes = 1, ylen, xlen ;
		clay:_DeflateLevel = 1 ;

	short cfvo(depth, lat, lon) ;
		cfvo:long_name = "coarse fragments by volume" ;
		cfvo:units = "fraction" ;
		cfvo:_FillValue = -32768s ;
		cfvo:missing_value = -32768s ;
		cfvo:actual_range = 100.f, -100.f ;
		cfvo:valid_range = 0s, 1000s ;
		cfvo:scale_factor = 0.001f ;
		cfvo:_Storage = "chunked" ;
		cfvo:_Shuffle = "true" ;
		cfvo:_ChunkSizes = 1, ylen, xlen ;
		cfvo:_DeflateLevel = 1 ;

	short soc(depth, lat, lon) ;
		soc:long_name = "Soil organic carbon content by mass" ;
		soc:units = "fraction" ;
		soc:_FillValue = -32768s ;
		soc:missing_value = -32768s ;
		soc:actual_range = 100.f, -100.f ;
		soc:valid_range = 0s, 10000s ;
		soc:scale_factor = 0.0001f ;
		soc:_Storage = "chunked" ;
		soc:_Shuffle = "true" ;
		soc:_ChunkSizes = 1, ylen, xlen ;
		soc:_DeflateLevel = 1 ;

	float Tsat(depth, lat, lon) ;
		Tsat:long_name = "soil porosity (Theta-sat)" ;
		Tsat:units = "fraction" ;
		Tsat:_FillValue = -9999.f ;
		Tsat:missing_value = -9999.f ;
		Tsat:actual_range = 0.f, 1.f ;
		Tsat:_Storage = "chunked" ;
		Tsat:_ChunkSizes = 1, ylen, xlen ;
		Tsat:_DeflateLevel = 1 ;

	float whc(depth, lat, lon) ;
		whc:long_name = "water holding capacity defined as T33-T1500, reduced for coarse fragment volume" ;
		whc:units = "mm cm-1" ;
		whc:_FillValue = -9999.f ;
		whc:missing_value = -9999.f ;
		whc:actual_range = 0.f, 1000.f ;
		whc:_Storage = "chunked" ;
		whc:_ChunkSizes = 1, ylen, xlen ;
		whc:_DeflateLevel = 1 ;

	float Ksat(depth, lat, lon) ;
		Ksat:long_name = "saturated hydraulic conductivity" ;
		Ksat:units = "mm h-1" ;
		Ksat:_FillValue = -9999.f ;
		Ksat:missing_value = -9999.f ;
		Ksat:actual_range = 100.f, -100.f ;
		Ksat:_Storage = "chunked" ;
		Ksat:_ChunkSizes = 1, ylen, xlen ;

// global attributes:
		:Conventions = "CF-1.11" ;
		:title = "Primary and derived soil properties" ;
		:data_sources = "SoilGrids 250m (2020)" ;
		:node_offset = 1 ;

}
